----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:28:19 04/23/2020 
-- Design Name: 
-- Module Name:    bin_to_bcd - Behavioral 
-- Project Name: 	 Ultrasonic_range_detector
-- Target Devices: CoolRunner-II CPLD starter board
-- Tool versions: 
-- Description: 	 Module for retyping distance from std_logic_vector to binary decimal code
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity bin_to_bcd is
port(
		in
end bin_to_bcd;

architecture Behavioral of bin_to_bcd is

begin


end Behavioral;

